LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY AESKey IS
    PORT (
        KeyO   : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"000102030405060708090a0b0c0d0e0f";
        KeyR1  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"d6aa74fdd2af72fadaa678f1d6ab76fe";
        KeyR2  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"b692cf0b643dbdf1be9bc5006830b3fe";
        KeyR3  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"b6ff744ed2c2c9bf6c590cbf0469bf41";
        KeyR4  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"47f7f7bc95353e03f96c32bcfd058dfd";
        KeyR5  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"3caaa3e8a99f9deb50f3af57adf622aa";
        KeyR6  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"5e390f7df7a69296a7553dc10aa31f6b";
        KeyR7  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"14f9701ae35fe28c440adf4d4ea9c026";
        KeyR8  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"47438735a41c65b9e016baf4aebf7ad2";
        KeyR9  : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"549932d1f08557681093ed9cbe2c974e";
        KeyR10 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0) := x"13111d7fe3944a17f307a78b4d2b30c5"
    );
END AESKey;

ARCHITECTURE Behavioral OF AESKey IS

BEGIN
END Behavioral;